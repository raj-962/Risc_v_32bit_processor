module instruction_mem(
    input clk,
    input rst,
    input [31:0] read_addr,
    output reg [31:0] instruction_out
);

    reg [31:0] I_Mem[0:63]; // 64 instructions max
 integer i;
    // Combinational read
    always @(*) begin
        instruction_out = I_Mem[read_addr >> 2]; // Word-aligned access
    end

    // Initialize instructions
    initial begin
       
        // Clear memory
        for (i = 0; i < 64; i = i + 1) begin
            I_Mem[i] = 32'h00000000;
        end

  I_Mem[0] = 32'b0000000000000000000000000000000 ;       // no operation
        I_Mem[1] = 32'b0000000_11001_10000_000_01101_0110011;    // add x13, x16, x25
        I_Mem[2] = 32'b0100000_00011_01000_000_00101_0110011;     // sub x5, x8, x3
        I_Mem[3] = 32'b0000000_00011_00010_111_00001_0110011;    // and x1, x2, x3
        I_Mem[4] = 32'b0000000_00101_00011_110_00100_0110011;    // or x4, x3, x5
        I_Mem[5] = 32'b0000000_00101_00011_100_00100_0110011;    // xor x4, x3, x5
	    I_Mem[6] = 32'b0000000_00101_00011_001_00100_0110011;    // sll x4, x3, x5
        I_Mem[7] = 32'b0000000_00101_00011_101_00100_0110011;    // srl x4, x3, x5
        I_Mem[8] = 32'b0100000_00010_00011_101_00101_0110011;    //sra x5, x3, x2
        I_Mem[9] = 32'b0000000_00010_00011_010_00101_0110011;    //slt x5, x3, x2 
        // I-type
        I_Mem[10]  = 32'b000000000010_10101_000_10110_0010011;     // addi x22, x21, 2
        I_Mem[11]  = 32'b000000000011_01000_110_01001_0010011;     // ori x9, x8, 3 
	    I_Mem[12] = 32'b000000000100_01000_110_01001_0010011;     // xori x9, x8, 4
	    I_Mem[13] = 32'b000000000101_00010_111_00001_0010011;     // andi x1, x2, 5
	    I_Mem[14] = 32'b000000000110_00011_001_00100_0010011;    // slli x4, x3, 6
	    I_Mem[15] = 32'b000000000111_00011_101_00100_0010011;    // srli x4, x3, 7 
	    I_Mem[16] = 32'b000000001000_00011_101_00101_0010011;    //srai x5, x3, 8
	    I_Mem[17] = 32'b000000001001_00011_010_00101_0010011;    //slti x5, x3, 9  
        // L-type
	    I_Mem[18]=  32'b000000000101_00011_000_01001_0000011;     // lb x9, 5(x3)
	    I_Mem[19] = 32'b000000000011_00011_001_01001_0000011;    // lh x9, 3(x3)
        I_Mem[20]= 32'b000000001111_00010_010_01000_0000011;    // lw x8, 15(x2) 
        // S-type
        I_Mem[21] =  32'b0000000_01111_00011_000_01000_0100011;     // sb x15, 8(x3), x3 = 12
	    I_Mem[22] =  32'b0000000_01110_00110_001_01010_0100011;     // sh x14, 10(x6), x6 = 44
	    I_Mem[23] = 32'b0000000_01110_00110_010_01100_0100011;     // sw x14, 12(x6), x6 = 44     
	//B-type    
	    I_Mem[24] = 32'b0_000000_01001_01001_000_0110_0_1100011;     // beq x9, x9, 12, (PC + 12 if x9 = x9 
	    I_Mem[25] = 32'b0_000000_01001_01001_001_0111_0_1100011;     //bne x9, x9, 14,(PC + 14 if x9 != x9)
	// U-type
        I_Mem[26] =  32'b00000000000000101000_00011_0110111;     // lui x3, 40
        I_Mem[27] =  32'b0000000000000010100_00101_0010111;     // auipc x5, 20 (rd = PC + (imm << 12))
	// J-type
	    I_Mem[28] = 32'b0_00000000_0_0000010100_00001_1101111;         // jal x1, 20

    end

endmodule